module nand1(input  wire a, b,
             output wire y);
  assign y = ~(a & b);
endmodule